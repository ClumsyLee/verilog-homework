module data_whiting(
    output reg [9:0] tx_data,
    output reg tx_valid,
    output reg rx_ready,
    input [9:0] rx_data,
    input rx_status,
    input next_rx_ready,
    input clk,
    input reset_n
);



endmodule
