module serial_transceiver(dout, din, clk);

output dout;
input din, clk;



endmodule
