module framing_encoding(
    output reg framing_encoding_out,
    output reg framing_encoding_out_valid,
    input [7:0] phr_psdu_in,
    input phr_psdu_in_valid,
    input clk,
    input reset_n
);



endmodule
